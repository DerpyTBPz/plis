library verilog;
use verilog.vl_types.all;
entity testbench is
    generic(
        CLK_PERIOD      : integer := 125
    );
end testbench;
