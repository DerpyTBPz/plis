library verilog;
use verilog.vl_types.all;
entity testbench2 is
    generic(
        CLK_PERIOD      : integer := 125
    );
end testbench2;
